
package OOP_tb_pkg;

    `include "ALU_reference_model.sv"
    `include "alu_trans.sv"
    `include "generator.sv"
    `include "driver.sv"
    `include "monitor_inputs.sv"
    `include "monitor_outputs.sv"
    `include "scoreboard.sv"
    `include "coverg.sv"
    `include "env.sv"

endpackage