package alu_pkg;
import uvm_pkg::*;


`include "uvm_macros.svh"
`include "ALU_reference_model.sv"
`include "seq_item.sv"
`include "random_sequence.sv"
`include "sequencer.sv"
`include "driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"
`include "coverage.sv"
`include "agent.sv"
`include "environment.sv"
`include "test.sv"  


endpackage